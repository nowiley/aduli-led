`timescale 1ns / 1ps
`include "mem/xilinx_single_port_ram_read_first.v"
`include "calibration/id_shower.sv"
`default_nettype none

module cal_fsm
endmodule

`default_nettype wire